module main

fn main(){
	s := "Hello World!"
	x := 1
	d := 2.2

	println("Printing variables")
	println("Printing text: ${s}")
	println("Printing integer: ${x}")
	println("Printing decimal: ${d}")
}
